library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.STD_LOGIC_arith.all;
use ieee.STD_LOGIC_unsigned.all;

entity memory_m is
-- memory_m port 
	port(  
		memory_write: in STD_LOGIC;
		clk: in STD_LOGIC;
		data_in : in STD_LOGIC_VECTOR(15 downto 0);
		address : in STD_LOGIC_VECTOR(15 downto 0);
		data_out : out STD_LOGIC_VECTOR(15 downto 0)
	);
end memory_m;

architecture behavioral of memory_m is


-- creating array 
type mem_array is array(0 to 511) of STD_LOGIC_VECTOR(15 downto 0);

begin

memory_m: process(data_in, memory_write, clk)
variable control_memory : mem_array:=(

-- 16 bits:
-- 0-6 = opcode
-- 7-9 = destanation address 
-- 10-12 = source A
-- 13-15 = source B

		-- 0
		x"0004", -- 0
		x"0006", -- 1
		x"0242", -- 2
		x"0B02", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"ABCD", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 1
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 2
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 3
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 4
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 5
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 6
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 7
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 8
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 9
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- A
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- B
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- C
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- D
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- E
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- F
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 0
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 1
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 2
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 3
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 4
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 5
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 6
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 7
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 8
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- 9
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- A
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- B
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- C
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- D
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- E
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000", -- F

		-- F
		x"0000", -- 0
		x"0000", -- 1
		x"0000", -- 2
		x"0000", -- 3
		x"0000", -- 4
		x"0000", -- 5
		x"0000", -- 6
		x"0000", -- 7
		x"0000", -- 8
		x"0000", -- 9
		x"0000", -- A
		x"0000", -- B
		x"0000", -- C
		x"0000", -- D
		x"0000", -- E
		x"0000"  -- F

	);

	variable int_addr : integer;
	variable cut_addr: STD_LOGIC_VECTOR(8 downto 0);
	variable array_output: STD_LOGIC_VECTOR(15 downto 0);


	begin 
		if (rising_edge(clk)) then
		
			cut_addr := address(8 downto 0);
			int_addr := conv_integer(cut_addr);

			if(memory_write = '0') then
			
				array_output := control_memory(int_addr);
				data_out <= array_output(15 downto 0);

			elsif (memory_write = '1') then 
			
				control_memory(int_addr) := data_in;

			else
			end if;
		end if;
	end process;
end behavioral;
